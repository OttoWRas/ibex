
package aespim_pkg;



endpackage : aespim_pkg